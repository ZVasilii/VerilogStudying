module tick(input clk, output clk_1);
    assign clk_1 = clk;
endmodule
